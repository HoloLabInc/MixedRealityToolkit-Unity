<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>Class ParabolaLineDataProvider
   | Mixed Reality Toolkit Documentation </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="Class ParabolaLineDataProvider
   | Mixed Reality Toolkit Documentation ">
    <meta name="generator" content="docfx 2.48.0.0">
    
    <link rel="shortcut icon" href=".././Documentation/Images/favicon.ico">
    <link rel="stylesheet" href="../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../styles/docfx.css">
    <link rel="stylesheet" href="../styles/main.css">
    <meta property="docfx:navrel" content="../toc.html">
    <meta property="docfx:tocrel" content="toc.html">
    
    <meta property="docfx:rel" content="../">
    
    <!-- Global site tag (gtag.js) - Google Analytics -->
    <script async="" src="https://www.googletagmanager.com/gtag/js?id=UA-177859076-1"></script>
    <script>
    window.dataLayer = window.dataLayer || [];
    function gtag(){dataLayer.push(arguments);}
    gtag('js', new Date());
  
    gtag('config', 'UA-177859076-1');
    </script>
  </head>
  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              
              <a class="navbar-brand" href="../index.html">
                <img id="logo" class="svg" src=".././Documentation/Images/mrt_logo_icon.png" alt="">
              </a>
            </div>
          
          <div class="version-dropdown" id="versionDropdown">
           </div>
         
          <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div class="container body-content">
        
        <div id="search-results">
          <div class="search-list"></div>
          <div class="sr-items">
            <p><i class="glyphicon glyphicon-refresh index-loading"></i></p>
          </div>
          <ul id="pagination"></ul>
        </div>
      </div>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider">
  
  
  <h1 id="Microsoft_MixedReality_Toolkit_Utilities_ParabolaLineDataProvider" data-uid="Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider" class="text-break">Class ParabolaLineDataProvider
  </h1>
  <div class="markdown level0 summary"><p sourcefile="../../obj/api/Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.yml" sourcestartlinenumber="2">Base Parabola line data provider.</p>
</div>
  <div class="markdown level0 conceptual"></div>
  <div class="inheritance">
    <h5>Inheritance</h5>
    <div class="level0"><a class="xref" href="https://docs.microsoft.com/dotnet/api/system.object">Object</a></div>
    <div class="level1"><a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html">BaseMixedRealityLineDataProvider</a></div>
    <div class="level2"><span class="xref">ParabolaLineDataProvider</span></div>
      <div class="level3"><a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.ParabolaConstrainedLineDataProvider.html">ParabolaConstrainedLineDataProvider</a></div>
      <div class="level3"><a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.ParabolaPhysicalLineDataProvider.html">ParabolaPhysicalLineDataProvider</a></div>
  </div>
  <div class="inheritedMembers">
    <h5>Inherited Members</h5>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_LineStartClamp">BaseMixedRealityLineDataProvider.LineStartClamp</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_LineEndClamp">BaseMixedRealityLineDataProvider.LineEndClamp</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_LineTransform">BaseMixedRealityLineDataProvider.LineTransform</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_Loops">BaseMixedRealityLineDataProvider.Loops</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_TransformMode">BaseMixedRealityLineDataProvider.TransformMode</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_RotationMode">BaseMixedRealityLineDataProvider.RotationMode</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_FlipUpVector">BaseMixedRealityLineDataProvider.FlipUpVector</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_OriginOffset">BaseMixedRealityLineDataProvider.OriginOffset</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_ManualUpVectorBlend">BaseMixedRealityLineDataProvider.ManualUpVectorBlend</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_ManualUpVectors">BaseMixedRealityLineDataProvider.ManualUpVectors</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_VelocitySearchRange">BaseMixedRealityLineDataProvider.VelocitySearchRange</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_Distorters">BaseMixedRealityLineDataProvider.Distorters</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_DistortionEnabled">BaseMixedRealityLineDataProvider.DistortionEnabled</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_DistortionMode">BaseMixedRealityLineDataProvider.DistortionMode</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_DistortionStrength">BaseMixedRealityLineDataProvider.DistortionStrength</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_UniformDistortionStrength">BaseMixedRealityLineDataProvider.UniformDistortionStrength</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_FirstPoint">BaseMixedRealityLineDataProvider.FirstPoint</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_LastPoint">BaseMixedRealityLineDataProvider.LastPoint</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_UnClampedWorldLength">BaseMixedRealityLineDataProvider.UnClampedWorldLength</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_PointCount">BaseMixedRealityLineDataProvider.PointCount</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_SetPointInternal_System_Int32_Vector3_">BaseMixedRealityLineDataProvider.SetPointInternal(Int32, Vector3)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetPointInternal_System_Single_">BaseMixedRealityLineDataProvider.GetPointInternal(Single)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetPointInternal_System_Int32_">BaseMixedRealityLineDataProvider.GetPointInternal(Int32)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_UnclampedWorldLengthSearchSteps">BaseMixedRealityLineDataProvider.UnclampedWorldLengthSearchSteps</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_OnEnable">BaseMixedRealityLineDataProvider.OnEnable()</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_LateUpdate">BaseMixedRealityLineDataProvider.LateUpdate()</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetNormalizedLengthFromWorldLength_System_Single_System_Int32_">BaseMixedRealityLineDataProvider.GetNormalizedLengthFromWorldLength(Single, Int32)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetVelocity_System_Single_">BaseMixedRealityLineDataProvider.GetVelocity(Single)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetRotation_System_Single_Microsoft_MixedReality_Toolkit_LineRotationMode_">BaseMixedRealityLineDataProvider.GetRotation(Single, LineRotationMode)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetRotation_System_Int32_Microsoft_MixedReality_Toolkit_LineRotationMode_">BaseMixedRealityLineDataProvider.GetRotation(Int32, LineRotationMode)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetPoint_System_Single_">BaseMixedRealityLineDataProvider.GetPoint(Single)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetUnClampedPoint_System_Single_">BaseMixedRealityLineDataProvider.GetUnClampedPoint(Single)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetPoint_System_Int32_">BaseMixedRealityLineDataProvider.GetPoint(Int32)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_SetPoint_System_Int32_Vector3_">BaseMixedRealityLineDataProvider.SetPoint(Int32, Vector3)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetClosestPoint_Vector3_System_Int32_System_Int32_">BaseMixedRealityLineDataProvider.GetClosestPoint(Vector3, Int32, Int32)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetNormalizedLengthFromWorldPos_Vector3_System_Int32_System_Int32_">BaseMixedRealityLineDataProvider.GetNormalizedLengthFromWorldPos(Vector3, Int32, Int32)</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_UpdateMatrix">BaseMixedRealityLineDataProvider.UpdateMatrix()</a>
    </div>
    <div>
      <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_DrawUnselectedGizmosPreview">BaseMixedRealityLineDataProvider.DrawUnselectedGizmosPreview()</a>
    </div>
  </div>
  <h6><strong>Namespace</strong>: <a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.html">Microsoft.MixedReality.Toolkit.Utilities</a></h6>
  <h6><strong>Assembly</strong>: cs.temp.dll.dll</h6>
  <h5 id="Microsoft_MixedReality_Toolkit_Utilities_ParabolaLineDataProvider_syntax">Syntax</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">public abstract class ParabolaLineDataProvider : BaseMixedRealityLineDataProvider</code></pre>
  </div>
  <h3 id="properties">Properties
  </h3>
  
  
  <a id="Microsoft_MixedReality_Toolkit_Utilities_ParabolaLineDataProvider_StartPoint_" data-uid="Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.StartPoint*"></a>
  <h4 id="Microsoft_MixedReality_Toolkit_Utilities_ParabolaLineDataProvider_StartPoint" data-uid="Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.StartPoint">StartPoint</h4>
  <div class="markdown level1 summary"><p sourcefile="../../obj/api/Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.yml" sourcestartlinenumber="2">The Starting point of this line.</p>
</div>
  <div class="markdown level1 conceptual"></div>
  <h5 class="decalaration">Declaration</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">public MixedRealityPose StartPoint { get; }</code></pre>
  </div>
  <h5 class="propertyValue">Property Value</h5>
  <table class="table table-bordered table-striped table-condensed">
    <thead>
      <tr>
        <th>Type</th>
        <th>Description</th>
      </tr>
    </thead>
    <tbody>
      <tr>
        <td><a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.MixedRealityPose.html">MixedRealityPose</a></td>
        <td></td>
      </tr>
    </tbody>
  </table>
  <h5 id="Microsoft_MixedReality_Toolkit_Utilities_ParabolaLineDataProvider_StartPoint_remarks">Remarks</h5>
  <div class="markdown level1 remarks"><p sourcefile="../../obj/api/Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.yml" sourcestartlinenumber="1">Always located at this <a href="https://docs.unity3d.com/ScriptReference/GameObject.html">GameObject</a>'s <a href="https://docs.unity3d.com/ScriptReference/Transform-position.html">Transform.position</a></p>
</div>
  <h3 id="methods">Methods
  </h3>
  
  
  <a id="Microsoft_MixedReality_Toolkit_Utilities_ParabolaLineDataProvider_GetUnClampedWorldLengthInternal_" data-uid="Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.GetUnClampedWorldLengthInternal*"></a>
  <h4 id="Microsoft_MixedReality_Toolkit_Utilities_ParabolaLineDataProvider_GetUnClampedWorldLengthInternal" data-uid="Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.GetUnClampedWorldLengthInternal">GetUnClampedWorldLengthInternal()</h4>
  <div class="markdown level1 summary"><p sourcefile="../../obj/api/Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.yml" sourcestartlinenumber="2">Get the UnClamped world length of the line</p>
</div>
  <div class="markdown level1 conceptual"></div>
  <h5 class="decalaration">Declaration</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">protected override float GetUnClampedWorldLengthInternal()</code></pre>
  </div>
  <h5 class="returns">Returns</h5>
  <table class="table table-bordered table-striped table-condensed">
    <thead>
      <tr>
        <th>Type</th>
        <th>Description</th>
      </tr>
    </thead>
    <tbody>
      <tr>
        <td><a class="xref" href="https://docs.microsoft.com/dotnet/api/system.single">Single</a></td>
        <td></td>
      </tr>
    </tbody>
  </table>
  <h5 class="overrides">Overrides</h5>
  <div><a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetUnClampedWorldLengthInternal">BaseMixedRealityLineDataProvider.GetUnClampedWorldLengthInternal()</a></div>
  
  
  <a id="Microsoft_MixedReality_Toolkit_Utilities_ParabolaLineDataProvider_GetUpVectorInternal_" data-uid="Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.GetUpVectorInternal*"></a>
  <h4 id="Microsoft_MixedReality_Toolkit_Utilities_ParabolaLineDataProvider_GetUpVectorInternal_System_Single_" data-uid="Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.GetUpVectorInternal(System.Single)">GetUpVectorInternal(Single)</h4>
  <div class="markdown level1 summary"><p sourcefile="../../obj/api/Microsoft.MixedReality.Toolkit.Utilities.ParabolaLineDataProvider.yml" sourcestartlinenumber="2">Gets the up vector at a normalized length along line (used for rotation)</p>
</div>
  <div class="markdown level1 conceptual"></div>
  <h5 class="decalaration">Declaration</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">protected override Vector3 GetUpVectorInternal(float normalizedLength)</code></pre>
  </div>
  <h5 class="parameters">Parameters</h5>
  <table class="table table-bordered table-striped table-condensed">
    <thead>
      <tr>
        <th>Type</th>
        <th>Name</th>
        <th>Description</th>
      </tr>
    </thead>
    <tbody>
      <tr>
        <td><a class="xref" href="https://docs.microsoft.com/dotnet/api/system.single">Single</a></td>
        <td><span class="parametername">normalizedLength</span></td>
        <td></td>
      </tr>
    </tbody>
  </table>
  <h5 class="returns">Returns</h5>
  <table class="table table-bordered table-striped table-condensed">
    <thead>
      <tr>
        <th>Type</th>
        <th>Description</th>
      </tr>
    </thead>
    <tbody>
      <tr>
        <td><span class="xref">Vector3</span></td>
        <td></td>
      </tr>
    </tbody>
  </table>
  <h5 class="overrides">Overrides</h5>
  <div><a class="xref" href="Microsoft.MixedReality.Toolkit.Utilities.BaseMixedRealityLineDataProvider.html#Microsoft_MixedReality_Toolkit_Utilities_BaseMixedRealityLineDataProvider_GetUpVectorInternal_System_Single_">BaseMixedRealityLineDataProvider.GetUpVectorInternal(Single)</a></div>
</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
              <!-- <p><a class="back-to-top" href="#top">Back to top</a><p> -->
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            
            <span>Generated by <strong>DocFX</strong></span>
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../styles/docfx.js"></script>
    <script type="text/javascript" src="../styles/main.js"></script>
  </body>
</html>
