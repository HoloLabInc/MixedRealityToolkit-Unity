a   �  a   v     0  �  �    *  ]  r  \  p  y  �  �  �  �  �  �  �  �  �     v   FileAndType�     �{"baseDir":"D:/a/1/s/scripts/docs","file":"../../Documentation.ja/README_NearMenu.md","type":"article","sourceDir":"../../","destinationDir":"./"}   0  OriginalFileAndType�   �  �{"baseDir":"D:/a/1/s/scripts/docs","file":"../../Documentation.ja/README_NearMenu.md","type":"article","sourceDir":"../../","destinationDir":"./"}   �  Key5     +~/../../Documentation.ja/README_NearMenu.md   *  LocalPathFromRoot3   ]  )../../Documentation.ja/README_NearMenu.md   r  LinkToFilesA   \  �  �  H  |  �    P  �  �    `  �  �    L   �  B~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom2.pngI   H  ?~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Grab.png4   |  *~/../../Documentation.ja/README_Sliders.mdN   �  D~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Structure.png:     0~/../../Documentation.ja/README_BoundsControl.mdL   P  B~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom1.pngD   �  :~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu.pngL   �  B~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom0.png3     )~/../../Documentation.ja/README_Button.mdM   `  C~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Examples.png@   �  6~/../../Documentation.ja/README_ManipulationHandler.mdL   �  B~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom3.png3     )~/../../Documentation.ja/README_Solver.md=   \  3~/../../Documentation.ja/README_ObjectCollection.md   p  
LinkToUids	   y     �  FileLinkSources  �  �{"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom2.png":[{"Target":"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom2.png","LineNumber":0}],"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Grab.png":[{"Target":"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Grab.png","LineNumber":0}],"~/../../Documentation.ja/README_Sliders.md":[{"Target":"~/../../Documentation.ja/README_Sliders.md","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":69}],"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Structure.png":[{"Target":"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Structure.png","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":41}],"~/../../Documentation.ja/README_BoundsControl.md":[{"Target":"~/../../Documentation.ja/README_BoundsControl.md","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":68}],"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom1.png":[{"Target":"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom1.png","LineNumber":0}],"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu.png":[{"Target":"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu.png","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":3}],"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom0.png":[{"Target":"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom0.png","LineNumber":0}],"~/../../Documentation.ja/README_Button.md":[{"Target":"~/../../Documentation.ja/README_Button.md","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":36},{"Target":"~/../../Documentation.ja/README_Button.md","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":67}],"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Examples.png":[{"Target":"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Examples.png","LineNumber":0}],"~/../../Documentation.ja/README_ManipulationHandler.md":[{"Target":"~/../../Documentation.ja/README_ManipulationHandler.md","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":38},{"Target":"~/../../Documentation.ja/README_ManipulationHandler.md","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":71}],"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom3.png":[{"Target":"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom3.png","LineNumber":0}],"~/../../Documentation.ja/README_Solver.md":[{"Target":"~/../../Documentation.ja/README_Solver.md","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":39},{"Target":"~/../../Documentation.ja/README_Solver.md","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":72}],"~/../../Documentation.ja/README_ObjectCollection.md":[{"Target":"~/../../Documentation.ja/README_ObjectCollection.md","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":37},{"Target":"~/../../Documentation.ja/README_ObjectCollection.md","SourceFile":"../../Documentation.ja/README_NearMenu.md","LineNumber":70}]}   �  UidLinkSources   �  {}   �  Uids   �  []   �  ManifestProperties�   �  �{"rawTitle":"<h1 id=\"near-menu\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"1\">Near menu</h1>"}   �  DocumentType	   �   �6  IJ  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","conceptual":"\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"3\"><img src=\"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu.png\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"3\" alt=\"Near Menu\"></p>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"5\">Near Menu is a UX control which provides a collection of buttons or other UI components. It is floating around the user's body and easily accessible anytime. Since it is loosely coupled with the user, it does not disturb the user's interaction with the target content. The user can use the 'Pin' button to world-lock/unlock the menu. The menu can be grabbed and placed at a specific position.</p>\n<h2 id=\"interaction-behavior\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"7\">Interaction behavior</h2>\n<ul sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"9\">\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"9\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"9\">Tag-along</strong>: The menu follows you and stays within 30-60cm range from the user for the near interactions.</li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"10\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"10\">Pin</strong>: Using the 'Pin' button, the menu can be world-locked and released.</li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"11\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"11\">Grab and move</strong>: The menu is always grabbable and movable. Regardless of the previous state, the menu will be pinned(world-locked) when grabbed and released. There are visual cues for the grabbable area. They are revealed on hand proximity.</li>\n</ul>\n<img src=\"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Grab.png\">\n<h2 id=\"prefabs\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"15\">Prefabs</h2>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"17\">Near Menu prefabs are designed to demonstrate how to use MRTK's various components to build menus for near interactions.</p>\n<ul sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"19\">\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"19\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"19\">NearMenu2x4.prefab</strong></li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"20\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"20\">NearMenu3x1.prefab</strong></li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"21\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"21\">NearMenu3x2.prefab</strong></li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"22\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"22\">NearMenu3x3.prefab</strong></li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"23\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"23\">NearMenu4x1.prefab</strong></li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"24\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"24\">NearMenu4x2.prefab</strong></li>\n</ul>\n<h2 id=\"example-scene\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"26\">Example scene</h2>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"28\">You can find examples of Near Menu prefabs in the <code sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"28\">NearMenuExamples</code> scene.</p>\n<img src=\"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Examples.png\">\n<h2 id=\"structure\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"32\">Structure</h2>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"34\">Near Menu prefabs are made with following MRTK components.</p>\n<ul sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"36\">\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"36\"><a href=\"~/../../Documentation.ja/README_Button.md\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"36\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"36\">PressableButtonHoloLens2</strong></a> prefab</li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"37\"><a href=\"~/../../Documentation.ja/README_ObjectCollection.md\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"37\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"37\">Grid Object Collection</strong></a>: Multiple button layout in grid</li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"38\"><a href=\"~/../../Documentation.ja/README_ManipulationHandler.md\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"38\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"38\">Manipulation Handler</strong></a>: Grab and move the menu</li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"39\"><a href=\"~/../../Documentation.ja/README_Solver.md\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"39\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"39\">RadialView Solver</strong></a>: Follow Me(tag-along) behavior</li>\n</ul>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"41\"><img src=\"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Structure.png\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"41\" alt=\"Near Menu Prefab\"></p>\n<h2 id=\"how-to-customize\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"43\">How to customize</h2>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"45\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"45\">1. Add/Remove Buttons</strong></p>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"47\">Under <code sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"47\">ButtonCollection</code> object, add or remove buttons.<br>\n<img src=\"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom0.png\" width=\"450\"></p>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"50\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"50\">2. Update the Grid Object Collection</strong></p>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"52\">Click <code sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"52\">Update Collection</code> button in the Inspector of the <code sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"52\">ButtonCollection</code> object. It will update the grid layout.<br>\n<img src=\"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom1.png\"></p>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"55\">You can configure the number of rows using <code sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"55\">Rows</code> property of the Grid Object Collection.<br>\n<img src=\"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom2.png\"></p>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"58\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"58\">3. Adjust the backplate size</strong></p>\n<p sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"60\">Adjust the size of the <code sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"60\">Quad</code> under <code sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"60\">Backplate</code> object. The width and height of the backplate should be <code sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"60\">0.032 * [Number of the buttons + 1]</code>. For example, if you have 3 x 2 buttons, the width of the backplate is <code sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"60\">0.032 * 4</code> and the height is <code sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"60\">0.032 * 3</code>. You can directly put this expression into the Unity's field.<br>\n<img src=\"~/../../Documentation/Images/NearMenu/MRTK_UX_NearMenu_Custom3.png\" width=\"450\"></p>\n<ul sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"63\">\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"63\">Default size of the HoloLens 2 button is 3.2x3.2 cm (0.032m)</li>\n</ul>\n<h2 id=\"see-also\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"65\">See also</h2>\n<ul sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"67\">\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"67\"><a href=\"~/../../Documentation.ja/README_Button.md\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"67\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"67\">Buttons</strong></a></li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"68\"><a href=\"~/../../Documentation.ja/README_BoundsControl.md\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"68\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"68\">Bounds Control</strong></a></li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"69\"><a href=\"~/../../Documentation.ja/README_Sliders.md\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"69\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"69\">Slider</strong></a></li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"70\"><a href=\"~/../../Documentation.ja/README_ObjectCollection.md\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"70\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"70\">Grid Object Collection</strong></a></li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"71\"><a href=\"~/../../Documentation.ja/README_ManipulationHandler.md\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"71\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"71\">Manipulation Handler</strong></a></li>\n<li sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"72\"><a href=\"~/../../Documentation.ja/README_Solver.md\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"72\"><strong sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"72\">RadialView Solver</strong></a></li>\n</ul>\n","type":"Conceptual","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"Documentation.ja/README_NearMenu.md","branch":"mrtk_documentation_ja","repo":"https://github.com/HoloLabInc/MixedRealityToolkit-Unity"},"startLine":0,"endLine":0,"isExternal":false},"path":"../../Documentation.ja/README_NearMenu.md","documentation":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"Documentation.ja/README_NearMenu.md","branch":"mrtk_documentation_ja","repo":"https://github.com/HoloLabInc/MixedRealityToolkit-Unity"},"startLine":0,"endLine":0,"isExternal":false},"_enableSearch":true,"_docfxVersion":"2.48.0.0","_disableNavbar":false,"_appLogoPath":"./Documentation/Images/mrt_logo_icon.png","_gitContribute":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","repo":"https://github.com/Microsoft/MixedRealityToolkit-Unity","branch":"mrtk_development"},"_appFaviconPath":"./Documentation/Images/favicon.ico","_appTitle":"Mixed Reality Toolkit Documentation","_systemKeys":{"$type":"System.String[], mscorlib","$values":["conceptual","type","source","path","documentation","title","rawTitle","wordCount"]},"rawTitle":"<h1 id=\"near-menu\" sourcefile=\"../../Documentation.ja/README_NearMenu.md\" sourcestartlinenumber=\"1\">Near menu</h1>","title":"Near menu"}�   �J  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","IsUserDefinedTitle":false,"XrefSpec":null}	   �J   